module _16_to_23_decoder(d,q); // this module is 16 to 23 decorder module
input [15:0] d; // define 16 bits input d
output reg [22:0] q; // define 23 bits output q and 23 bits reg q

always @ (d) // Calculate the next state through the case statement
begin // begin - end means { }
	case(d) 
	16'h0100 : q = 23'b0000000000_0000000000_001;
	16'h0101 : q = 23'b0000000000_0000000000_010;
	16'h0102 : q = 23'b0000000000_0000000000_100;
	16'h0103 : q = 23'b0000000000_0000000001_000;
	16'h0104 : q = 23'b0000000000_0000000010_000;
	16'h0105 : q = 23'b0000000000_0000000100_000;
	16'h0106 : q = 23'b0000000000_0000001000_000;
	16'h0107 : q = 23'b0000000000_0000010000_000;
	16'h0108 : q = 23'b0000000000_0000100000_000;
	16'h0109 : q = 23'b0000000000_0001000000_000;
	16'h0110 : q = 23'b0000000000_0010000000_000;
	16'h0111 : q = 23'b0000000000_0100000000_000;
	16'h0112 : q = 23'b0000000000_1000000000_000;
	16'h0113 : q = 23'b0000000001_0000000000_000;
	16'h0114 : q = 23'b0000000010_0000000000_000;
	16'h0115 : q = 23'b0000000100_0000000000_000;
	16'h0116 : q = 23'b0000001000_0000000000_000;
	16'h0117 : q = 23'b0000010000_0000000000_000;
	16'h0118 : q = 23'b0000100000_0000000000_000;
	16'h0119 : q = 23'b0001000000_0000000000_000;
	16'h0120 : q = 23'b0010000000_0000000000_000;
	16'h0121 : q = 23'b0100000000_0000000000_000;
	16'h0122 : q = 23'b1000000000_0000000000_000;
	default : q = 23'hx; // To prevent the problem of latch
	endcase // end of case
end
endmodule // end of module